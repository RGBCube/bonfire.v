module bonfire

// hello_world prints "Hello, world!" to the console.
pub fn hello_world() {
	println('Hello, world!')
}
